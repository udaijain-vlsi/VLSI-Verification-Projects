module fifo (
input clk,
input rst,
input wr_en,      
input rd_en,      
input [7:0] data_in,
output reg [7:0] data_out,
output full,
output empty,
output reg led        
);
reg [7:0] memory [0:7];   
reg [2:0] wr_ptr, rd_ptr;
reg [3:0] count;
assign full  = (count == 8);
assign empty = (count == 0);
always @(posedge clk or posedge rst) begin
if (rst) begin
wr_ptr <= 0;
rd_ptr <= 0;
count  <= 0;
led    <= 0;
end
else begin
if (wr_en && !full) begin
memory[wr_ptr] <= data_in;
wr_ptr <= wr_ptr + 1;
count  <= count + 1;
end
if (rd_en && !empty) begin
data_out <= memory[rd_ptr];
rd_ptr <= rd_ptr + 1;
count  <= count - 1;
end
led <= full;
end
end
endmodule
